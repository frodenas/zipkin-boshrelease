CREATE KEYSPACE IF NOT EXISTS "Zipkin" WITH replication = {'class': 'SimpleStrategy', 'replication_factor': 1};

CREATE TABLE IF NOT EXISTS "Zipkin"."Traces" (
    key blob,
    column1 blob,
    value blob,
    PRIMARY KEY (key, column1)
) WITH CLUSTERING ORDER BY (column1 ASC)
    AND COMPACT STORAGE
    AND compaction = {'min_threshold': '4', 'class': 'org.apache.cassandra.db.compaction.SizeTieredCompactionStrategy', 'max_threshold': '32'};

CREATE TABLE IF NOT EXISTS "Zipkin"."SpanNames" (
    key blob,
    column1 blob,
    value blob,
    PRIMARY KEY (key, column1)
) WITH CLUSTERING ORDER BY (column1 ASC)
    AND COMPACT STORAGE
    AND compaction = {'min_threshold': '4', 'class': 'org.apache.cassandra.db.compaction.SizeTieredCompactionStrategy', 'max_threshold': '32'};

CREATE TABLE IF NOT EXISTS "Zipkin"."ServiceNames" (
    key blob,
    column1 blob,
    value blob,
    PRIMARY KEY (key, column1)
) WITH CLUSTERING ORDER BY (column1 ASC)
    AND COMPACT STORAGE
    AND compaction = {'min_threshold': '4', 'class': 'org.apache.cassandra.db.compaction.SizeTieredCompactionStrategy', 'max_threshold': '32'};

CREATE TABLE IF NOT EXISTS "Zipkin"."ServiceNameIndex" (
    key blob,
    column1 bigint,
    value blob,
    PRIMARY KEY (key, column1)
) WITH CLUSTERING ORDER BY (column1 ASC)
    AND COMPACT STORAGE
    AND compaction = {'min_threshold': '4', 'class': 'org.apache.cassandra.db.compaction.SizeTieredCompactionStrategy', 'max_threshold': '32'};

CREATE TABLE IF NOT EXISTS "Zipkin"."ServiceSpanNameIndex" (
    key blob,
    column1 bigint,
    value blob,
    PRIMARY KEY (key, column1)
) WITH CLUSTERING ORDER BY (column1 ASC)
    AND COMPACT STORAGE
    AND compaction = {'min_threshold': '4', 'class': 'org.apache.cassandra.db.compaction.SizeTieredCompactionStrategy', 'max_threshold': '32'};

CREATE TABLE IF NOT EXISTS "Zipkin"."AnnotationsIndex" (
    key blob,
    column1 bigint,
    value blob,
    PRIMARY KEY (key, column1)
) WITH CLUSTERING ORDER BY (column1 ASC)
    AND COMPACT STORAGE
    AND compaction = {'min_threshold': '4', 'class': 'org.apache.cassandra.db.compaction.SizeTieredCompactionStrategy', 'max_threshold': '32'};

CREATE TABLE IF NOT EXISTS "Zipkin"."Dependencies" (
    key blob,
    column1 bigint,
    value blob,
    PRIMARY KEY (key, column1)
) WITH CLUSTERING ORDER BY (column1 ASC)
    AND COMPACT STORAGE
    AND compaction = {'min_threshold': '4', 'class': 'org.apache.cassandra.db.compaction.SizeTieredCompactionStrategy', 'max_threshold': '32'};

CREATE TABLE IF NOT EXISTS "Zipkin"."DurationIndex" (
    key blob,
    column1 bigint,
    value blob,
    PRIMARY KEY (key, column1)
) WITH CLUSTERING ORDER BY (column1 ASC)
    AND COMPACT STORAGE
    AND compaction = {'min_threshold': '4', 'class': 'org.apache.cassandra.db.compaction.SizeTieredCompactionStrategy', 'max_threshold': '32'};

CREATE TABLE IF NOT EXISTS "Zipkin"."TopAnnotations" (
    key blob,
    column1 bigint,
    value blob,
    PRIMARY KEY (key, column1)
) WITH CLUSTERING ORDER BY (column1 ASC)
    AND COMPACT STORAGE
    AND compaction = {'min_threshold': '4', 'class': 'org.apache.cassandra.db.compaction.SizeTieredCompactionStrategy', 'max_threshold': '32'};
